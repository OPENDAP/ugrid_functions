netcdf hex {
dimensions:
	time = 3 ;
	faces = 8 ;
	nodes = 9 ;
	three = 3 ;
variables:
	int fvcom_mesh ;
		fvcom_mesh:face_node_connectivity = "fnca" ;
		fvcom_mesh:standard_name = "mesh_topology" ;
		fvcom_mesh:dimension = 2 ;
		fvcom_mesh:node_coordinates = "X Y" ;
	float X(nodes) ;
		X:grid = "element" ;
		X:grid_location = "node" ;
	float Y(nodes) ;
		Y:grid = "element" ;
		Y:grid_location = "node" ;
	int fnca(three, faces) ;
		fnca:start_index = 1 ;
		fnca:standard_name = "face_node_connectivity" ;
	float oneDnodedata(nodes) ;
		oneDnodedata:coordinates = "Y X" ;
		oneDnodedata:mesh = "fvcom_mesh" ;
		oneDnodedata:location = "node" ;
	float twoDnodedata(time, nodes) ;
		oneDnodedata:coordinates = "Y X" ;
		oneDnodedata:mesh = "fvcom_mesh" ;
		oneDnodedata:location = "node" ;
	float celldata(faces) ;
		celldata:mesh = "fvcom_mesh" ;
		celldata:location = "face" ;
	float bogusMeshRef(nodes) ;
		bogusMeshRef:coordinates = "Y X" ;
		bogusMeshRef:mesh = "bogus" ;
		bogusMeshRef:location = "node" ;
data:

 fvcom_mesh = 666;
 
 X = -1.0, 0.0, 1.0, 1.5,  1.0,  0.0, -1.0, -1.5, 0.0 ;

 Y =  1.0, 1.5, 1.0, 0.0, -1.0, -1.5, -1.0,  0.0, 0.0 ;

 fnca =
  1, 2, 3, 4, 5, 6, 7, 8,
  2, 3, 4, 5, 6, 7, 8, 1,
  9, 9, 9, 9, 9, 9, 9, 9;

 oneDnodedata = 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9;
 
 twoDnodedata = 
  0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9,
  1.1, 1.2, 1.3, 1.4, 1.5, 1.6, 1.7, 1.8, 1.9,
  2.1, 2.2, 2.3, 2.4, 2.5, 2.6, 2.7, 2.8, 2.9;

 celldata = 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8 ;
 
 bogusMeshRef = 0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 0.7, 0.8, 0.9;

}
